/*
*  File            :   pwm.svh
*  Autor           :   Vlasov D.V.
*  Data            :   2019.07.11
*  Language        :   SystemVerilog
*  Description     :   This is PWM module header file
*  Copyright(c)    :   2019 Vlasov D.V.
*/

`ifndef PWM_DEFS
`define PWM_DEFS
    parameter PWM_C_R = 'h0;
`endif
