/*
*  File            :   gpio.svh
*  Autor           :   Vlasov D.V.
*  Data            :   2019.07.11
*  Language        :   SystemVerilog
*  Description     :   This is GPIO module header file
*  Copyright(c)    :   2019 Vlasov D.V.
*/

`ifndef GPIO_DEFS
`define GPIO_DEFS
    parameter GPIO_GPI_R = 'h0;
    parameter GPIO_GPO_R = 'h4;
    parameter GPIO_GPD_R = 'h8;
`endif
