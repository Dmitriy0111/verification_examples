`ifndef TEST_PARAM_PKG__SVH
`define TEST_PARAM_PKG__SVH

package test_param_pkg;

    parameter DW = 587;

endpackage : test_param_pkg

`endif // TEST_PARAM_PKG__SVH
